library verilog;
use verilog.vl_types.all;
entity c3_vlg_vec_tst is
end c3_vlg_vec_tst;
