library verilog;
use verilog.vl_types.all;
entity c2_vlg_vec_tst is
end c2_vlg_vec_tst;
